/////////////////////////////////////////////////////////////////////////
//                                                                     //
//   Modulename :  sys_defs.svh                                        //
//                                                                     //
//  Description :  This file has the macro-defines for macros used in  //
//                 the pipeline design.                                //
//                                                                     //
/////////////////////////////////////////////////////////////////////////

`ifndef __SYS_DEFS_SVH__
`define __SYS_DEFS_SVH__

// NOTE: moved this into sys_defs.svh, don't add to any other files
// have all files `include "sys_defs.svh" from now on (why weren't we doing this before?)
`timescale 1ns/100ps

// Synthesis testing definition for parameterized modules tested at multiple sizes
// see lab 6 CAM for example usage
`ifdef SYNTH_TEST
`define INSTANCE(mod) mod``_svsim
`else
`define INSTANCE(mod) mod
`endif

//////////////////////////////////////////////
//
// Memory/testbench attribute definitions
//
//////////////////////////////////////////////

// NOTE: the CLOCK_PERIOD definition has been moved to the Makefile

// cache mode removes the byte-level interface from memory, so it always returns a double word
// the original processor won't work with this defined
// so your new processor will have to account for our changes to mem
`define CACHE_MODE // MUST BE DEFINED FOR FINAL PROCESSOR

// you are not allowed to change this definition for your final processor
`define MEM_LATENCY_IN_CYCLES (100.0/`CLOCK_PERIOD+0.49999)
// the 0.49999 is to force ceiling(100/period). The default behavior for
// float to integer conversion is rounding to nearest

// the original p3 definition - can be useful for temporarily testing non-memory functionality
// `define MEM_LATENCY_IN_CYCLES 0


`define NUM_MEM_TAGS 15

`define MEM_SIZE_IN_BYTES (64*1024)
`define MEM_64BIT_LINES   (`MEM_SIZE_IN_BYTES/8)

typedef union packed {
    logic [7:0][7:0]  byte_level;
    logic [3:0][15:0] half_level;
    logic [1:0][31:0] word_level;
} EXAMPLE_CACHE_BLOCK;

`ifndef CACHE_MODE
typedef enum logic [1:0] {
	BYTE = 2'h0,
	HALF = 2'h1,
	WORD = 2'h2,
	DOUBLE = 2'h3
} MEM_SIZE;
`endif


//////////////////////////////////////////////
// Exception codes
// This mostly follows the RISC-V Privileged spec
// except a few add-ons for our infrastructure
// The majority of them won't be used, but it's
// good to know what they are
//////////////////////////////////////////////

typedef enum logic [3:0] {
	INST_ADDR_MISALIGN  = 4'h0,
	INST_ACCESS_FAULT   = 4'h1,
	ILLEGAL_INST        = 4'h2,
	BREAKPOINT          = 4'h3,
	LOAD_ADDR_MISALIGN  = 4'h4,
	LOAD_ACCESS_FAULT   = 4'h5,
	STORE_ADDR_MISALIGN = 4'h6,
	STORE_ACCESS_FAULT  = 4'h7,
	ECALL_U_MODE        = 4'h8,
	ECALL_S_MODE        = 4'h9,
	NO_ERROR            = 4'ha, //a reserved code that we modified for our purpose
	ECALL_M_MODE        = 4'hb,
	INST_PAGE_FAULT     = 4'hc,
	LOAD_PAGE_FAULT     = 4'hd,
	HALTED_ON_WFI       = 4'he, //another reserved code that we used
	STORE_PAGE_FAULT    = 4'hf
} EXCEPTION_CODE;

//////////////////////////////////////////////
//
// Datapath control signals
//
//////////////////////////////////////////////

// ALU opA input mux selects
typedef enum logic [1:0] {
	OPA_IS_RS1  = 2'h0,
	OPA_IS_NPC  = 2'h1,
	OPA_IS_PC   = 2'h2,
	OPA_IS_ZERO = 2'h3
} ALU_OPA_SELECT;

// ALU opB input mux selects
typedef enum logic [3:0] {
	OPB_IS_RS2    = 4'h0,
	OPB_IS_I_IMM  = 4'h1,
	OPB_IS_S_IMM  = 4'h2,
	OPB_IS_B_IMM  = 4'h3,
	OPB_IS_U_IMM  = 4'h4,
	OPB_IS_J_IMM  = 4'h5
} ALU_OPB_SELECT;

// Destination register select
typedef enum logic [1:0] {
	DEST_RD = 2'h0,
	DEST_NONE  = 2'h1
} DEST_REG_SEL;

// ALU function code input
// probably want to leave these alone
typedef enum logic [4:0] {
	ALU_ADD     = 5'h00,
	ALU_SUB     = 5'h01,
	ALU_SLT     = 5'h02,
	ALU_SLTU    = 5'h03,
	ALU_AND     = 5'h04,
	ALU_OR      = 5'h05,
	ALU_XOR     = 5'h06,
	ALU_SLL     = 5'h07,
	ALU_SRL     = 5'h08,
	ALU_SRA     = 5'h09,
	ALU_MUL     = 5'h0a,
	ALU_MULH    = 5'h0b,
	ALU_MULHSU  = 5'h0c,
	ALU_MULHU   = 5'h0d,
	ALU_DIV     = 5'h0e,
	ALU_DIVU    = 5'h0f,
	ALU_REM     = 5'h10,
	ALU_REMU    = 5'h11
} ALU_FUNC;

//////////////////////////////////////////////
//
// Assorted things it is not wise to change
//
//////////////////////////////////////////////

// actually, you might have to change this if you change VERILOG_CLOCK_PERIOD
// JK you don't ^^^
`define SD #1

// the RISCV register file zero register, any read of this register always
// returns a zero value, and any write to this register is thrown away
`define ZERO_REG 5'd0

// Memory bus commands control signals
typedef enum logic [1:0] {
	BUS_NONE     = 2'h0,
	BUS_LOAD     = 2'h1,
	BUS_STORE    = 2'h2
} BUS_COMMAND;

`ifndef CACHE_MODE
typedef enum logic [1:0] {
	BYTE = 2'h0,
	HALF = 2'h1,
	WORD = 2'h2,
	DOUBLE = 2'h3
} MEM_SIZE;
`endif

// useful boolean single-bit definitions
`define FALSE  1'h0
`define TRUE  1'h1

// RISCV ISA SPEC
`define XLEN 32
typedef union packed {
	logic [31:0] inst;
	struct packed {
		logic [6:0] funct7;
		logic [4:0] rs2;
		logic [4:0] rs1;
		logic [2:0] funct3;
		logic [4:0] rd;
		logic [6:0] opcode;
	} r; //register to register instructions
	struct packed {
		logic [11:0] imm;
		logic [4:0]  rs1; //base
		logic [2:0]  funct3;
		logic [4:0]  rd;  //dest
		logic [6:0]  opcode;
	} i; //immediate or load instructions
	struct packed {
		logic [6:0] off; //offset[11:5] for calculating address
		logic [4:0] rs2; //source
		logic [4:0] rs1; //base
		logic [2:0] funct3;
		logic [4:0] set; //offset[4:0] for calculating address
		logic [6:0] opcode;
	} s; //store instructions
	struct packed {
		logic       of;  //offset[12]
		logic [5:0] s;   //offset[10:5]
		logic [4:0] rs2; //source 2
		logic [4:0] rs1; //source 1
		logic [2:0] funct3;
		logic [3:0] et;  //offset[4:1]
		logic       f;   //offset[11]
		logic [6:0] opcode;
	} b; //branch instructions
	struct packed {
		logic [19:0] imm;
		logic [4:0]  rd;
		logic [6:0]  opcode;
	} u; //upper immediate instructions
	struct packed {
		logic       of; //offset[20]
		logic [9:0] et; //offset[10:1]
		logic       s;  //offset[11]
		logic [7:0] f;	//offset[19:12]
		logic [4:0] rd; //dest
		logic [6:0] opcode;
	} j;  //jump instructions
`ifdef ATOMIC_EXT
	struct packed {
		logic [4:0] funct5;
		logic       aq;
		logic       rl;
		logic [4:0] rs2;
		logic [4:0] rs1;
		logic [2:0] funct3;
		logic [4:0] rd;
		logic [6:0] opcode;
	} a; //atomic instructions
`endif
`ifdef SYSTEM_EXT
	struct packed {
		logic [11:0] csr;
		logic [4:0]  rs1;
		logic [2:0]  funct3;
		logic [4:0]  rd;
		logic [6:0]  opcode;
	} sys; //system call instructions
`endif

} INST; //instruction typedef, this should cover all types of instructions

//
// Basic NOP instruction.  Allows pipline registers to clearly be reset with
// an instruction that does nothing instead of Zero which is really an ADDI x0, x0, 0
//
`define NOP 32'h00000013

//////////////////////////////////////////////
//
// IF Packets:
// Data that is exchanged between the IF and the ID stages
//
//////////////////////////////////////////////

typedef struct packed {
	logic valid; // If low, the data in this struct is garbage
    INST  inst;  // fetched instruction out
	logic [`XLEN-1:0] NPC; // PC + 4
	logic [`XLEN-1:0] PC;  // PC
} IF_ID_PACKET;

//////////////////////////////////////////////
//
// ID Packets:
// Data that is exchanged from ID to EX stage
//
//////////////////////////////////////////////

typedef struct packed {
	logic [`XLEN-1:0] NPC; // PC + 4
	logic [`XLEN-1:0] PC;  // PC

	logic [`XLEN-1:0] rs1_value; // reg A value
	logic [`XLEN-1:0] rs2_value; // reg B value
	
	ALU_OPA_SELECT opa_select; // ALU opa mux select (ALU_OPA_xxx *)
	ALU_OPB_SELECT opb_select; // ALU opb mux select (ALU_OPB_xxx *)
	INST inst;                 // instruction
	
	logic [4:0] dest_reg_idx;  // destination (writeback) register index
	ALU_FUNC    alu_func;      // ALU function select (ALU_xxx *)
	logic       rd_mem;        // does inst read memory?
	logic       wr_mem;        // does inst write memory?
	logic       cond_branch;   // is inst a conditional branch?
	logic       uncond_branch; // is inst an unconditional branch?
	logic       halt;          // is this a halt?
	logic       illegal;       // is this instruction illegal?
	logic       csr_op;        // is this a CSR operation? (we only used this as a cheap way to get return code)
	logic       valid;         // is inst a valid instruction to be counted for CPI calculations?
} ID_EX_PACKET;

typedef struct packed {
	logic [`XLEN-1:0] alu_result;  // alu_result
	logic [`XLEN-1:0] NPC;         // pc + 4
	logic             take_branch; // is this a taken branch?
	// pass-through from decode stage
	logic [`XLEN-1:0] rs2_value;
	logic             rd_mem, wr_mem;
	logic [4:0]       dest_reg_idx;
	logic             halt, illegal, csr_op, valid;
	logic [2:0]       mem_size; // byte, half-word or word
} EX_MEM_PACKET;


//////////////////////////////////////////////
//
// NEW Project4 Packets:
// Packets used in Project4
//
//////////////////////////////////////////////

`define INST_LEN 32
`define REG_LEN $clog2(`INST_LEN)

`define ROB_LEN 8
`define RS_LEN 8
`define SUPERSCALER_LEN 1
`define MAP_TABLE_LEN 32
`define BTB_LEN 32


// flags for cdb write through
typedef enum logic [1:0] {TAGTAG, TAGCDB, CDBTAG, CDBCDB} FLAG;

// indicate which channel in ex
typedef enum logic [2:0] {ALU, MULT, BR, LD, ST} CHANNEL;

// packet of tag
typedef struct packed {
	logic [$clog2(`ROB_LEN)-1:0] tag;   //ROB entry number
	logic 						 valid; //valid bit (e.g. tag = 0 && valid = 1 => ROB#0, tag = 0 && valid = 0 => tag is empty)
} TAG_PACKET;

//////////////////////////////////////////////
//
// ID_packet:
// Data from decoder to RS in dispatch stage
//
//////////////////////////////////////////////

typedef struct packed {
	logic [`XLEN-1:0] NPC; // PC + 4
	logic [`XLEN-1:0] PC;  // PC

	logic [`XLEN-1:0] rs1_value; // reg A value
	logic [`XLEN-1:0] rs2_value; // reg B value
	
	ALU_OPA_SELECT opa_select; // ALU opa mux select (ALU_OPA_xxx *)
	ALU_OPB_SELECT opb_select; // ALU opb mux select (ALU_OPB_xxx *)
	INST inst;                 // instruction
	
	logic [4:0] dest_reg_idx;  // destination (writeback) register index
	ALU_FUNC    alu_func;      // ALU function select (ALU_xxx *)
	logic       rd_mem;        // does inst read memory?
	logic       wr_mem;        // does inst write memory?
	logic       cond_branch;   // is inst a conditional branch?
	logic       uncond_branch; // is inst an unconditional branch?
	logic       halt;          // is this a halt?
	logic       illegal;       // is this instruction illegal?
	logic       csr_op;        // is this a CSR operation? (we only used this as a cheap way to get return code)
	logic       valid;         // is inst a valid instruction to be counted for CPI calculations?
	CHANNEL     channel;
} ID_PACKET;

//////////////////////////////////////////////
//
// IS_packet:
// Data after D_S pipeline
//
//////////////////////////////////////////////

typedef struct packed {
	logic [`XLEN-1:0] NPC; // PC + 4
	logic [`XLEN-1:0] PC;  // PC

	logic [`XLEN-1:0] rs1_value; // reg A value
	logic [`XLEN-1:0] rs2_value; // reg B value
	
	ALU_OPA_SELECT opa_select; // ALU opa mux select (ALU_OPA_xxx *)
	ALU_OPB_SELECT opb_select; // ALU opb mux select (ALU_OPB_xxx *)
	INST inst;                 // instruction
	
	logic [$clog2(`ROB_LEN)-1:0] dest_reg_idx;  // destination (writeback) register rob entry number
	ALU_FUNC    alu_func;      // ALU function select (ALU_xxx *)
	logic       rd_mem;        // does inst read memory?
	logic       wr_mem;        // does inst write memory?
	logic       cond_branch;   // is inst a conditional branch?
	logic       uncond_branch; // is inst an unconditional branch?
	logic       halt;          // is this a halt?
	logic       illegal;       // is this instruction illegal?
	logic       csr_op;        // is this a CSR operation? (we only used this as a cheap way to get return code)
	logic       valid;         // is inst a valid instruction to be counted for CPI calculations?
} IS_PACKET;

//////////////////////////////////////////////
//
// MT2RS_PACKET:
// Data from Map Table to RS
//
//////////////////////////////////////////////

typedef struct packed {
	TAG_PACKET rs1_tag;
	TAG_PACKET rs2_tag;
	logic rs1_ready;
	logic rs2_ready;
} MT2RS_PACKET;

//////////////////////////////////////////////
//
// RS2MT_PACKET:
// Data from RS to Map Table
//
//////////////////////////////////////////////

typedef struct packed {
	logic [`REG_LEN-1:0] rs1_idx;
	logic [`REG_LEN-1:0] rs2_idx;
	logic [`REG_LEN-1:0] dest_reg_idx;
	TAG_PACKET dest_reg_tag;
} RS2MT_PACKET;

//////////////////////////////////////////////
//
// ROB2MT_PACKET:
// Data from ROB to Map Table
//
//////////////////////////////////////////////

typedef struct packed {
	logic retire;
	logic [$clog2(`ROB_LEN)-1:0] head_idx;
	logic squash;
} ROB2MT_PACKET;

//////////////////////////////////////////////
//
// CDB_PACKET:
// Data broadcasted from CDB
//
//////////////////////////////////////////////

typedef struct packed {
	TAG_PACKET reg_tag;
	logic [`XLEN-1:0] reg_value;
} CDB_PACKET;

//////////////////////////////////////////////
//
// ROB2RS_PACKET:
// Data from ROB to RS
//
//////////////////////////////////////////////

typedef struct packed {
	logic [$clog2(`ROB_LEN)-1:0] rob_entry;
	logic [$clog2(`ROB_LEN)-1:0] rob_head_idx;
	logic [`XLEN-1:0] rs1_value;
	logic [`XLEN-1:0] rs2_value;
	logic squash;
	//logic RS_enable;
} ROB2RS_PACKET;

//////////////////////////////////////////////
//
// RS2ROB_PACKET:
// Data from RS to ROB
//
//////////////////////////////////////////////

typedef struct packed {
	logic valid;
	logic [$clog2(`ROB_LEN)-1:0] rs1_idx;
	logic [$clog2(`ROB_LEN)-1:0] rs2_idx;
} RS2ROB_PACKET;

//////////////////////////////////////////////
//
// ROB_entry_PACKET:
// Data from ROB_entry to ROB
//
//////////////////////////////////////////////

typedef struct packed {
	logic [$clog2(`ROB_LEN)-1:0] dest_reg_value;  //data
	logic [$clog2(`ROB_LEN)-1:0] dest_reg_idx;    //address
	logic                        valid;
} ROB_entry_PACKET;

typedef struct packed {
	logic [`XLEN-1:0] alu_result;  // alu_result
	logic [`XLEN-1:0] NPC;         // pc + 4
	logic             take_branch; // is this a taken branch?
	logic [4:0]       dest_reg_idx;
	logic [`XLEN-1:0] rs2_value;	//rs2_value
	logic 			  stru_hazard; //if there is a structural hazard

	logic       	  rd_mem;        // does inst read memory?
	logic       	  wr_mem;        // does inst write memory?
	logic       	  cond_branch;   // is inst a conditional branch?
	logic       	  uncond_branch; // is inst an unconditional branch?
	logic       	  halt;          // is this a halt?
	logic       	  illegal;       // is this instruction illegal?
	logic       	  csr_op;        // is this a CSR operation? (we only used this as a cheap way to get return code)
	logic       	  valid;         // is inst a valid instruction to be counted for CPI calculations?
	logic [2:0]       mem_size;

} EX_OUT_PACKET;

typedef struct packed {
	TAG_PACKET mispredict_rob_entry_idx;
} MISPREDICT_ROB_PACKET;


//////////////////////////////////////////////
//
// ROB_entry_PACKET:
// Data from ROB_entry to ROB
//
//////////////////////////////////////////////
typedef struct packed {
	logic [`XLEN-1:0]    dest_reg_value;
	logic [`REG_LEN-1:0] dest_reg_idx;
} ROB2REG_PACKET;


//////////////////////////////////////////////
//
// IF2BTB_PACKET:
// Data from IF/ID to BTB
//
//////////////////////////////////////////////

typedef struct packed {
	logic [`XLEN-1:0] inst;
	logic valid;
} IFID2BTB_PACKET;


//////////////////////////////////////////////
//
// FU2BTB_PACKET:
// Data from Brcond FU to BTB
//
//////////////////////////////////////////////

typedef struct packed {
	logic [`XLEN-1:0] inst;
	logic [`XLEN-1:0] target_pc;
	logic valid;
	logic taken;
} FU2BTB_PACKET;


//////////////////////////////////////////////
//
// BTB_PACKET:
// Data from BTB
//
//////////////////////////////////////////////

typedef struct packed {
	logic prediction; // 0 for not taken and 1 for taken
	logic valid;
	logic [`XLEN-1:0] target_pc;
} BTB_PACKET;

//////////////////////////////////////////////
//
// BTB_ENTRY:
// Data from BTB
//
//////////////////////////////////////////////

typedef struct packed {
	BTB_PREDICT state; // T WT WN N
	logic busy;
	logic [`XLEN-1:$clog2(`BTB_LEN)] tag;
	logic [`XLEN-1:0] target_pc;
} BTB_ENTRY;

typedef enum {TAKEN, WEAK_TAKEN, WEAK_NOTTAKE, NOTTAKE} BTB_PREDICT;

`endif // __SYS_DEFS_SVH__
